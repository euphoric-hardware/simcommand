logic [15:0] image [484];
assign image[0] = 'd0;
assign image[1] = 'd0;
assign image[2] = 'd0;
assign image[3] = 'd0;
assign image[4] = 'd0;
assign image[5] = 'd0;
assign image[6] = 'd0;
assign image[7] = 'd0;
assign image[8] = 'd0;
assign image[9] = 'd0;
assign image[10] = 'd500;
assign image[11] = 'd49;
assign image[12] = 'd36;
assign image[13] = 'd133;
assign image[14] = 'd0;
assign image[15] = 'd0;
assign image[16] = 'd0;
assign image[17] = 'd0;
assign image[18] = 'd0;
assign image[19] = 'd0;
assign image[20] = 'd0;
assign image[21] = 'd0;
assign image[22] = 'd0;
assign image[23] = 'd0;
assign image[24] = 'd0;
assign image[25] = 'd0;
assign image[26] = 'd0;
assign image[27] = 'd0;
assign image[28] = 'd0;
assign image[29] = 'd0;
assign image[30] = 'd0;
assign image[31] = 'd0;
assign image[32] = 'd221;
assign image[33] = 'd15;
assign image[34] = 'd9;
assign image[35] = 'd30;
assign image[36] = 'd500;
assign image[37] = 'd0;
assign image[38] = 'd0;
assign image[39] = 'd0;
assign image[40] = 'd0;
assign image[41] = 'd0;
assign image[42] = 'd0;
assign image[43] = 'd0;
assign image[44] = 'd0;
assign image[45] = 'd0;
assign image[46] = 'd0;
assign image[47] = 'd0;
assign image[48] = 'd0;
assign image[49] = 'd0;
assign image[50] = 'd0;
assign image[51] = 'd0;
assign image[52] = 'd0;
assign image[53] = 'd0;
assign image[54] = 'd500;
assign image[55] = 'd42;
assign image[56] = 'd12;
assign image[57] = 'd14;
assign image[58] = 'd117;
assign image[59] = 'd0;
assign image[60] = 'd0;
assign image[61] = 'd0;
assign image[62] = 'd0;
assign image[63] = 'd0;
assign image[64] = 'd0;
assign image[65] = 'd0;
assign image[66] = 'd0;
assign image[67] = 'd0;
assign image[68] = 'd0;
assign image[69] = 'd0;
assign image[70] = 'd0;
assign image[71] = 'd0;
assign image[72] = 'd0;
assign image[73] = 'd0;
assign image[74] = 'd0;
assign image[75] = 'd0;
assign image[76] = 'd0;
assign image[77] = 'd500;
assign image[78] = 'd18;
assign image[79] = 'd9;
assign image[80] = 'd31;
assign image[81] = 'd500;
assign image[82] = 'd0;
assign image[83] = 'd0;
assign image[84] = 'd0;
assign image[85] = 'd0;
assign image[86] = 'd0;
assign image[87] = 'd0;
assign image[88] = 'd0;
assign image[89] = 'd0;
assign image[90] = 'd0;
assign image[91] = 'd0;
assign image[92] = 'd0;
assign image[93] = 'd0;
assign image[94] = 'd0;
assign image[95] = 'd0;
assign image[96] = 'd0;
assign image[97] = 'd0;
assign image[98] = 'd0;
assign image[99] = 'd0;
assign image[100] = 'd22;
assign image[101] = 'd8;
assign image[102] = 'd15;
assign image[103] = 'd332;
assign image[104] = 'd0;
assign image[105] = 'd0;
assign image[106] = 'd0;
assign image[107] = 'd0;
assign image[108] = 'd0;
assign image[109] = 'd0;
assign image[110] = 'd0;
assign image[111] = 'd0;
assign image[112] = 'd0;
assign image[113] = 'd0;
assign image[114] = 'd0;
assign image[115] = 'd0;
assign image[116] = 'd0;
assign image[117] = 'd0;
assign image[118] = 'd0;
assign image[119] = 'd0;
assign image[120] = 'd0;
assign image[121] = 'd0;
assign image[122] = 'd36;
assign image[123] = 'd10;
assign image[124] = 'd10;
assign image[125] = 'd74;
assign image[126] = 'd0;
assign image[127] = 'd0;
assign image[128] = 'd0;
assign image[129] = 'd0;
assign image[130] = 'd0;
assign image[131] = 'd0;
assign image[132] = 'd0;
assign image[133] = 'd0;
assign image[134] = 'd0;
assign image[135] = 'd0;
assign image[136] = 'd0;
assign image[137] = 'd0;
assign image[138] = 'd0;
assign image[139] = 'd0;
assign image[140] = 'd0;
assign image[141] = 'd0;
assign image[142] = 'd0;
assign image[143] = 'd0;
assign image[144] = 'd30;
assign image[145] = 'd9;
assign image[146] = 'd10;
assign image[147] = 'd69;
assign image[148] = 'd0;
assign image[149] = 'd0;
assign image[150] = 'd0;
assign image[151] = 'd0;
assign image[152] = 'd0;
assign image[153] = 'd0;
assign image[154] = 'd0;
assign image[155] = 'd0;
assign image[156] = 'd0;
assign image[157] = 'd0;
assign image[158] = 'd0;
assign image[159] = 'd0;
assign image[160] = 'd0;
assign image[161] = 'd0;
assign image[162] = 'd0;
assign image[163] = 'd0;
assign image[164] = 'd0;
assign image[165] = 'd0;
assign image[166] = 'd34;
assign image[167] = 'd10;
assign image[168] = 'd9;
assign image[169] = 'd57;
assign image[170] = 'd0;
assign image[171] = 'd0;
assign image[172] = 'd0;
assign image[173] = 'd0;
assign image[174] = 'd0;
assign image[175] = 'd0;
assign image[176] = 'd0;
assign image[177] = 'd0;
assign image[178] = 'd0;
assign image[179] = 'd0;
assign image[180] = 'd0;
assign image[181] = 'd0;
assign image[182] = 'd0;
assign image[183] = 'd0;
assign image[184] = 'd0;
assign image[185] = 'd125;
assign image[186] = 'd47;
assign image[187] = 'd43;
assign image[188] = 'd17;
assign image[189] = 'd9;
assign image[190] = 'd9;
assign image[191] = 'd42;
assign image[192] = 'd0;
assign image[193] = 'd0;
assign image[194] = 'd0;
assign image[195] = 'd0;
assign image[196] = 'd0;
assign image[197] = 'd0;
assign image[198] = 'd0;
assign image[199] = 'd0;
assign image[200] = 'd0;
assign image[201] = 'd0;
assign image[202] = 'd0;
assign image[203] = 'd0;
assign image[204] = 'd500;
assign image[205] = 'd91;
assign image[206] = 'd25;
assign image[207] = 'd14;
assign image[208] = 'd11;
assign image[209] = 'd10;
assign image[210] = 'd9;
assign image[211] = 'd8;
assign image[212] = 'd8;
assign image[213] = 'd11;
assign image[214] = 'd15;
assign image[215] = 'd16;
assign image[216] = 'd36;
assign image[217] = 'd0;
assign image[218] = 'd0;
assign image[219] = 'd0;
assign image[220] = 'd0;
assign image[221] = 'd0;
assign image[222] = 'd0;
assign image[223] = 'd0;
assign image[224] = 'd500;
assign image[225] = 'd91;
assign image[226] = 'd16;
assign image[227] = 'd11;
assign image[228] = 'd9;
assign image[229] = 'd8;
assign image[230] = 'd8;
assign image[231] = 'd8;
assign image[232] = 'd8;
assign image[233] = 'd8;
assign image[234] = 'd8;
assign image[235] = 'd8;
assign image[236] = 'd8;
assign image[237] = 'd8;
assign image[238] = 'd10;
assign image[239] = 'd41;
assign image[240] = 'd0;
assign image[241] = 'd0;
assign image[242] = 'd0;
assign image[243] = 'd0;
assign image[244] = 'd0;
assign image[245] = 'd500;
assign image[246] = 'd50;
assign image[247] = 'd14;
assign image[248] = 'd8;
assign image[249] = 'd8;
assign image[250] = 'd8;
assign image[251] = 'd8;
assign image[252] = 'd8;
assign image[253] = 'd8;
assign image[254] = 'd8;
assign image[255] = 'd8;
assign image[256] = 'd10;
assign image[257] = 'd10;
assign image[258] = 'd11;
assign image[259] = 'd10;
assign image[260] = 'd13;
assign image[261] = 'd50;
assign image[262] = 'd0;
assign image[263] = 'd0;
assign image[264] = 'd0;
assign image[265] = 'd0;
assign image[266] = 'd0;
assign image[267] = 'd166;
assign image[268] = 'd15;
assign image[269] = 'd8;
assign image[270] = 'd8;
assign image[271] = 'd8;
assign image[272] = 'd8;
assign image[273] = 'd8;
assign image[274] = 'd8;
assign image[275] = 'd8;
assign image[276] = 'd8;
assign image[277] = 'd10;
assign image[278] = 'd38;
assign image[279] = 'd80;
assign image[280] = 'd91;
assign image[281] = 'd69;
assign image[282] = 'd166;
assign image[283] = 'd0;
assign image[284] = 'd0;
assign image[285] = 'd0;
assign image[286] = 'd0;
assign image[287] = 'd0;
assign image[288] = 'd0;
assign image[289] = 'd181;
assign image[290] = 'd15;
assign image[291] = 'd8;
assign image[292] = 'd8;
assign image[293] = 'd8;
assign image[294] = 'd8;
assign image[295] = 'd8;
assign image[296] = 'd8;
assign image[297] = 'd8;
assign image[298] = 'd9;
assign image[299] = 'd18;
assign image[300] = 'd221;
assign image[301] = 'd0;
assign image[302] = 'd0;
assign image[303] = 'd0;
assign image[304] = 'd0;
assign image[305] = 'd0;
assign image[306] = 'd0;
assign image[307] = 'd0;
assign image[308] = 'd0;
assign image[309] = 'd0;
assign image[310] = 'd0;
assign image[311] = 'd221;
assign image[312] = 'd16;
assign image[313] = 'd8;
assign image[314] = 'd8;
assign image[315] = 'd8;
assign image[316] = 'd8;
assign image[317] = 'd8;
assign image[318] = 'd8;
assign image[319] = 'd10;
assign image[320] = 'd17;
assign image[321] = 'd71;
assign image[322] = 'd0;
assign image[323] = 'd0;
assign image[324] = 'd0;
assign image[325] = 'd0;
assign image[326] = 'd0;
assign image[327] = 'd0;
assign image[328] = 'd0;
assign image[329] = 'd0;
assign image[330] = 'd0;
assign image[331] = 'd0;
assign image[332] = 'd0;
assign image[333] = 'd199;
assign image[334] = 'd16;
assign image[335] = 'd9;
assign image[336] = 'd8;
assign image[337] = 'd8;
assign image[338] = 'd9;
assign image[339] = 'd10;
assign image[340] = 'd16;
assign image[341] = 'd54;
assign image[342] = 'd500;
assign image[343] = 'd500;
assign image[344] = 'd0;
assign image[345] = 'd0;
assign image[346] = 'd0;
assign image[347] = 'd0;
assign image[348] = 'd0;
assign image[349] = 'd0;
assign image[350] = 'd0;
assign image[351] = 'd0;
assign image[352] = 'd0;
assign image[353] = 'd0;
assign image[354] = 'd0;
assign image[355] = 'd0;
assign image[356] = 'd74;
assign image[357] = 'd23;
assign image[358] = 'd17;
assign image[359] = 'd17;
assign image[360] = 'd28;
assign image[361] = 'd51;
assign image[362] = 'd332;
assign image[363] = 'd0;
assign image[364] = 'd0;
assign image[365] = 'd0;
assign image[366] = 'd0;
assign image[367] = 'd0;
assign image[368] = 'd0;
assign image[369] = 'd0;
assign image[370] = 'd0;
assign image[371] = 'd0;
assign image[372] = 'd0;
assign image[373] = 'd0;
assign image[374] = 'd0;
assign image[375] = 'd0;
assign image[376] = 'd0;
assign image[377] = 'd0;
assign image[378] = 'd0;
assign image[379] = 'd0;
assign image[380] = 'd0;
assign image[381] = 'd0;
assign image[382] = 'd0;
assign image[383] = 'd0;
assign image[384] = 'd0;
assign image[385] = 'd0;
assign image[386] = 'd0;
assign image[387] = 'd0;
assign image[388] = 'd0;
assign image[389] = 'd0;
assign image[390] = 'd0;
assign image[391] = 'd0;
assign image[392] = 'd0;
assign image[393] = 'd0;
assign image[394] = 'd0;
assign image[395] = 'd0;
assign image[396] = 'd0;
assign image[397] = 'd0;
assign image[398] = 'd0;
assign image[399] = 'd0;
assign image[400] = 'd0;
assign image[401] = 'd0;
assign image[402] = 'd0;
assign image[403] = 'd0;
assign image[404] = 'd0;
assign image[405] = 'd0;
assign image[406] = 'd0;
assign image[407] = 'd0;
assign image[408] = 'd0;
assign image[409] = 'd0;
assign image[410] = 'd0;
assign image[411] = 'd0;
assign image[412] = 'd0;
assign image[413] = 'd0;
assign image[414] = 'd0;
assign image[415] = 'd0;
assign image[416] = 'd0;
assign image[417] = 'd0;
assign image[418] = 'd0;
assign image[419] = 'd0;
assign image[420] = 'd0;
assign image[421] = 'd0;
assign image[422] = 'd0;
assign image[423] = 'd0;
assign image[424] = 'd0;
assign image[425] = 'd0;
assign image[426] = 'd0;
assign image[427] = 'd0;
assign image[428] = 'd0;
assign image[429] = 'd0;
assign image[430] = 'd0;
assign image[431] = 'd0;
assign image[432] = 'd0;
assign image[433] = 'd0;
assign image[434] = 'd0;
assign image[435] = 'd0;
assign image[436] = 'd0;
assign image[437] = 'd0;
assign image[438] = 'd0;
assign image[439] = 'd0;
assign image[440] = 'd0;
assign image[441] = 'd0;
assign image[442] = 'd0;
assign image[443] = 'd0;
assign image[444] = 'd0;
assign image[445] = 'd0;
assign image[446] = 'd0;
assign image[447] = 'd0;
assign image[448] = 'd0;
assign image[449] = 'd0;
assign image[450] = 'd0;
assign image[451] = 'd0;
assign image[452] = 'd0;
assign image[453] = 'd0;
assign image[454] = 'd0;
assign image[455] = 'd0;
assign image[456] = 'd0;
assign image[457] = 'd0;
assign image[458] = 'd0;
assign image[459] = 'd0;
assign image[460] = 'd0;
assign image[461] = 'd0;
assign image[462] = 'd0;
assign image[463] = 'd0;
assign image[464] = 'd0;
assign image[465] = 'd0;
assign image[466] = 'd0;
assign image[467] = 'd0;
assign image[468] = 'd0;
assign image[469] = 'd0;
assign image[470] = 'd0;
assign image[471] = 'd0;
assign image[472] = 'd0;
assign image[473] = 'd0;
assign image[474] = 'd0;
assign image[475] = 'd0;
assign image[476] = 'd0;
assign image[477] = 'd0;
assign image[478] = 'd0;
assign image[479] = 'd0;
assign image[480] = 'd0;
assign image[481] = 'd0;
assign image[482] = 'd0;
assign image[483] = 'd0;
