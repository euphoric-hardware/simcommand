logic [15:0] results [108];
assign results[0] = 'd23;
assign results[1] = 'd22;
assign results[2] = 'd21;
assign results[3] = 'd20;
assign results[4] = 'd31;
assign results[5] = 'd30;
assign results[6] = 'd29;
assign results[7] = 'd28;
assign results[8] = 'd27;
assign results[9] = 'd26;
assign results[10] = 'd25;
assign results[11] = 'd24;
assign results[12] = 'd39;
assign results[13] = 'd38;
assign results[14] = 'd37;
assign results[15] = 'd36;
assign results[16] = 'd35;
assign results[17] = 'd60;
assign results[18] = 'd42;
assign results[19] = 'd55;
assign results[20] = 'd51;
assign results[21] = 'd48;
assign results[22] = 'd63;
assign results[23] = 'd101;
assign results[24] = 'd100;
assign results[25] = 'd104;
assign results[26] = 'd114;
assign results[27] = 'd158;
assign results[28] = 'd164;
assign results[29] = 'd50;
assign results[30] = 'd58;
assign results[31] = 'd85;
assign results[32] = 'd82;
assign results[33] = 'd88;
assign results[34] = 'd85;
assign results[35] = 'd93;
assign results[36] = 'd88;
assign results[37] = 'd85;
assign results[38] = 'd93;
assign results[39] = 'd88;
assign results[40] = 'd85;
assign results[41] = 'd93;
assign results[42] = 'd88;
assign results[43] = 'd88;
assign results[44] = 'd85;
assign results[45] = 'd93;
assign results[46] = 'd85;
assign results[47] = 'd93;
assign results[48] = 'd85;
assign results[49] = 'd93;
assign results[50] = 'd88;
assign results[51] = 'd85;
assign results[52] = 'd93;
assign results[53] = 'd88;
assign results[54] = 'd85;
assign results[55] = 'd93;
assign results[56] = 'd88;
assign results[57] = 'd85;
assign results[58] = 'd93;
assign results[59] = 'd88;
assign results[60] = 'd85;
assign results[61] = 'd93;
assign results[62] = 'd88;
assign results[63] = 'd93;
assign results[64] = 'd88;
assign results[65] = 'd85;
assign results[66] = 'd93;
assign results[67] = 'd88;
assign results[68] = 'd85;
assign results[69] = 'd93;
assign results[70] = 'd88;
assign results[71] = 'd93;
assign results[72] = 'd85;
assign results[73] = 'd88;
assign results[74] = 'd85;
assign results[75] = 'd93;
assign results[76] = 'd88;
assign results[77] = 'd93;
assign results[78] = 'd85;
assign results[79] = 'd88;
assign results[80] = 'd85;
assign results[81] = 'd88;
assign results[82] = 'd85;
assign results[83] = 'd88;
assign results[84] = 'd20;
assign results[85] = 'd85;
assign results[86] = 'd93;
assign results[87] = 'd88;
assign results[88] = 'd20;
assign results[89] = 'd85;
assign results[90] = 'd93;
assign results[91] = 'd88;
assign results[92] = 'd20;
assign results[93] = 'd85;
assign results[94] = 'd93;
assign results[95] = 'd88;
assign results[96] = 'd20;
assign results[97] = 'd85;
assign results[98] = 'd93;
assign results[99] = 'd88;
assign results[100] = 'd20;
assign results[101] = 'd85;
assign results[102] = 'd93;
assign results[103] = 'd88;
assign results[104] = 'd93;
assign results[105] = 'd20;
assign results[106] = 'd85;
assign results[107] = 'd88;
